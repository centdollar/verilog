// Shift register
// Author: Vincent Michelini
// Description: intended to make a shift register with a lot of modular
// functionality and paramaterization to make this functionality possible
//
// TODO: first get a basic shift register made.


module shift_reg
#(

)
(

    input [7 : 0] din_i,


);
