// Author: Vincent Michelini
// Description: verilog code for the FILO register, this will act as a stack
//              in future uses of this. Due to this the write and read enable
//              will be called push and pop respectively


module filo_reg
#(
    parameter DEPTH = 8,
    parameter WIDTH = 8
)
(
    
);
